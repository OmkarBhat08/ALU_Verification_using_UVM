`define WIDTH 8
`define COMMAND_WIDTH 4
`define POW_2_N $clog2(`WIDTH)
