`define WIDTH 8
`define COMMAND_WIDTH 4
